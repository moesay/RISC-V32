parameter ALU_ADD = 4'h0;
parameter ALU_SUB = 4'h1;
parameter ALU_AND = 4'h2;
parameter ALU_OR = 4'h3;
parameter ALU_XOR = 4'h4;
parameter ALU_SLL = 4'h5;
parameter ALU_SRL = 4'h6;
parameter ALU_SRA = 4'h7;
parameter ALU_SLT = 4'h8;
parameter ALU_SLTU = 4'h9;
parameter ALU_A_PASSTHROUGH = 4'hA;
parameter ALU_B_PASSTHROUGH = 4'hB;

parameter ALU_NOP = 4'hF;


parameter IMM_NONE = 3'h0;
parameter IMM_I = 3'h1;
parameter IMM_S = 3'h2;
parameter IMM_B = 3'h3;
parameter IMM_U = 3'h4;
parameter IMM_J = 3'h5;
